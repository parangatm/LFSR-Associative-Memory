`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 11.05.2020 20:54:37
// Design Name: 
// Module Name: Enable_Signal_Decoder
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module Enable_Signal_Decoder(input [3:0]X,output reg[15:0]Y);

    always@(*)
        begin
            case(X)
            4'b0000: Y=16'b1000_0000_0000_0000;
            4'b0001: Y=16'b1100_0000_0000_0000;
            4'b0010: Y=16'b0110_0000_0000_0000;
            4'b0011: Y=16'b0011_0000_0000_0000;
            4'b0100: Y=16'b0010_1000_0000_0000;
            4'b0101: Y=16'b0000_1100_0000_0000;
            4'b0110: Y=16'b0000_0110_0000_0000;
            4'b0111: Y=16'b0110_0011_0000_0000;
            4'b1000: Y=16'b0000_1000_1000_0000;
            4'b1001: Y=16'b0000_0010_0100_0000;
            4'b1010: Y=16'b0000_0000_1010_0000;
            4'b1011: Y=16'b0000_1001_1001_0000;
            4'b1100: Y=16'b0000_0000_1101_1000;
            4'b1101: Y=16'b0110_0000_0000_1100;
            4'b1110: Y=16'b0000_0000_0000_0110;
            4'b1111: Y=16'b0000_0000_0010_1101;
            endcase
        end
endmodule
